module notgate(
	input in,
	output out
);
	
	assign out = ~in;
	
endmodule
