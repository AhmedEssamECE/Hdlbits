module andgate( 
    input a, 
    input b, 
    output out );

endmodule
